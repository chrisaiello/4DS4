// experiment1b.v

// Generated using ACDS version 12.0sp2 263 at 2016.01.28.19:10:43

`timescale 1 ps / 1 ps
module experiment1b (
		input  wire [3:0]  push_button_i_external_connection_export,       //       push_button_i_external_connection.export
		input  wire [16:0] switch_i_external_connection_export,            //            switch_i_external_connection.export
		output wire [17:0] led_red_o_external_connection_export,           //           led_red_o_external_connection.export
		input  wire        clk_50_i_in_reset_reset_n,                      //                       clk_50_i_in_reset.reset_n
		input  wire        clk_50_i_in_clk,                                //                             clk_50_i_in.clk
		output wire [8:0]  led_green_o_external_connection_export,         //         led_green_o_external_connection.export
		output wire [6:0]  seven_segment_n_o_0_external_connection_export, // seven_segment_n_o_0_external_connection.export
		inout  wire [15:0] sram_0_external_interface_DQ,                   //               sram_0_external_interface.DQ
		output wire [17:0] sram_0_external_interface_ADDR,                 //                                        .ADDR
		output wire        sram_0_external_interface_LB_N,                 //                                        .LB_N
		output wire        sram_0_external_interface_UB_N,                 //                                        .UB_N
		output wire        sram_0_external_interface_CE_N,                 //                                        .CE_N
		output wire        sram_0_external_interface_OE_N,                 //                                        .OE_N
		output wire        sram_0_external_interface_WE_N                  //                                        .WE_N
	);

	wire         cpu_0_instruction_master_waitrequest;                                                                            // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire  [20:0] cpu_0_instruction_master_address;                                                                                // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire         cpu_0_instruction_master_read;                                                                                   // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire  [31:0] cpu_0_instruction_master_readdata;                                                                               // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire         cpu_0_data_master_waitrequest;                                                                                   // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                                                                     // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire  [20:0] cpu_0_data_master_address;                                                                                       // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire         cpu_0_data_master_write;                                                                                         // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire         cpu_0_data_master_read;                                                                                          // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire  [31:0] cpu_0_data_master_readdata;                                                                                      // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                                                                                   // cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                                                                    // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                // cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                  // cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                               // cpu_0_jtag_debug_module_translator:av_chipselect -> cpu_0:jtag_debug_module_select
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                    // cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                 // cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                            // cpu_0_jtag_debug_module_translator:av_begintransfer -> cpu_0:jtag_debug_module_begintransfer
	wire         cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                              // cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                               // cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire  [15:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                               // sram_0_avalon_sram_slave_translator:av_writedata -> sram_0:writedata
	wire  [17:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                                 // sram_0_avalon_sram_slave_translator:av_address -> sram_0:address
	wire         sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                                   // sram_0_avalon_sram_slave_translator:av_write -> sram_0:write
	wire         sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                                    // sram_0_avalon_sram_slave_translator:av_read -> sram_0:read
	wire  [15:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                                // sram_0:readdata -> sram_0_avalon_sram_slave_translator:av_readdata
	wire         sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                           // sram_0:readdatavalid -> sram_0_avalon_sram_slave_translator:av_readdatavalid
	wire   [1:0] sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                              // sram_0_avalon_sram_slave_translator:av_byteenable -> sram_0:byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                        // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                          // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                            // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                         // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                              // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                               // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                           // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] switch_i_s1_translator_avalon_anti_slave_0_writedata;                                                            // SWITCH_I_s1_translator:av_writedata -> SWITCH_I:writedata
	wire   [1:0] switch_i_s1_translator_avalon_anti_slave_0_address;                                                              // SWITCH_I_s1_translator:av_address -> SWITCH_I:address
	wire         switch_i_s1_translator_avalon_anti_slave_0_chipselect;                                                           // SWITCH_I_s1_translator:av_chipselect -> SWITCH_I:chipselect
	wire         switch_i_s1_translator_avalon_anti_slave_0_write;                                                                // SWITCH_I_s1_translator:av_write -> SWITCH_I:write_n
	wire  [31:0] switch_i_s1_translator_avalon_anti_slave_0_readdata;                                                             // SWITCH_I:readdata -> SWITCH_I_s1_translator:av_readdata
	wire  [31:0] push_button_i_s1_translator_avalon_anti_slave_0_writedata;                                                       // PUSH_BUTTON_I_s1_translator:av_writedata -> PUSH_BUTTON_I:writedata
	wire   [1:0] push_button_i_s1_translator_avalon_anti_slave_0_address;                                                         // PUSH_BUTTON_I_s1_translator:av_address -> PUSH_BUTTON_I:address
	wire         push_button_i_s1_translator_avalon_anti_slave_0_chipselect;                                                      // PUSH_BUTTON_I_s1_translator:av_chipselect -> PUSH_BUTTON_I:chipselect
	wire         push_button_i_s1_translator_avalon_anti_slave_0_write;                                                           // PUSH_BUTTON_I_s1_translator:av_write -> PUSH_BUTTON_I:write_n
	wire  [31:0] push_button_i_s1_translator_avalon_anti_slave_0_readdata;                                                        // PUSH_BUTTON_I:readdata -> PUSH_BUTTON_I_s1_translator:av_readdata
	wire  [31:0] led_red_o_s1_translator_avalon_anti_slave_0_writedata;                                                           // LED_RED_O_s1_translator:av_writedata -> LED_RED_O:writedata
	wire   [1:0] led_red_o_s1_translator_avalon_anti_slave_0_address;                                                             // LED_RED_O_s1_translator:av_address -> LED_RED_O:address
	wire         led_red_o_s1_translator_avalon_anti_slave_0_chipselect;                                                          // LED_RED_O_s1_translator:av_chipselect -> LED_RED_O:chipselect
	wire         led_red_o_s1_translator_avalon_anti_slave_0_write;                                                               // LED_RED_O_s1_translator:av_write -> LED_RED_O:write_n
	wire  [31:0] led_red_o_s1_translator_avalon_anti_slave_0_readdata;                                                            // LED_RED_O:readdata -> LED_RED_O_s1_translator:av_readdata
	wire  [31:0] led_green_o_s1_translator_avalon_anti_slave_0_writedata;                                                         // LED_GREEN_O_s1_translator:av_writedata -> LED_GREEN_O:writedata
	wire   [1:0] led_green_o_s1_translator_avalon_anti_slave_0_address;                                                           // LED_GREEN_O_s1_translator:av_address -> LED_GREEN_O:address
	wire         led_green_o_s1_translator_avalon_anti_slave_0_chipselect;                                                        // LED_GREEN_O_s1_translator:av_chipselect -> LED_GREEN_O:chipselect
	wire         led_green_o_s1_translator_avalon_anti_slave_0_write;                                                             // LED_GREEN_O_s1_translator:av_write -> LED_GREEN_O:write_n
	wire  [31:0] led_green_o_s1_translator_avalon_anti_slave_0_readdata;                                                          // LED_GREEN_O:readdata -> LED_GREEN_O_s1_translator:av_readdata
	wire  [31:0] custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                              // custom_counter_component_0_avalon_slave_0_translator:av_writedata -> custom_counter_component_0:writedata
	wire   [1:0] custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                // custom_counter_component_0_avalon_slave_0_translator:av_address -> custom_counter_component_0:address
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                             // custom_counter_component_0_avalon_slave_0_translator:av_chipselect -> custom_counter_component_0:chipselect
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                  // custom_counter_component_0_avalon_slave_0_translator:av_write -> custom_counter_component_0:write
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                   // custom_counter_component_0_avalon_slave_0_translator:av_read -> custom_counter_component_0:read
	wire  [31:0] custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                               // custom_counter_component_0:readdata -> custom_counter_component_0_avalon_slave_0_translator:av_readdata
	wire  [31:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                             // custom_counter_component2_0_avalon_slave_0_translator:av_writedata -> custom_counter_component2_0:writedata
	wire   [1:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                               // custom_counter_component2_0_avalon_slave_0_translator:av_address -> custom_counter_component2_0:address
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                            // custom_counter_component2_0_avalon_slave_0_translator:av_chipselect -> custom_counter_component2_0:chipselect
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                 // custom_counter_component2_0_avalon_slave_0_translator:av_write -> custom_counter_component2_0:write
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                  // custom_counter_component2_0_avalon_slave_0_translator:av_read -> custom_counter_component2_0:read
	wire  [31:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // custom_counter_component2_0:readdata -> custom_counter_component2_0_avalon_slave_0_translator:av_readdata
	wire  [31:0] seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // SEVEN_SEGMENT_N_O_0_s1_translator:av_writedata -> SEVEN_SEGMENT_N_O_0:writedata
	wire   [1:0] seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_address;                                                   // SEVEN_SEGMENT_N_O_0_s1_translator:av_address -> SEVEN_SEGMENT_N_O_0:address
	wire         seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // SEVEN_SEGMENT_N_O_0_s1_translator:av_chipselect -> SEVEN_SEGMENT_N_O_0:chipselect
	wire         seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_write;                                                     // SEVEN_SEGMENT_N_O_0_s1_translator:av_write -> SEVEN_SEGMENT_N_O_0:write_n
	wire  [31:0] seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // SEVEN_SEGMENT_N_O_0:readdata -> SEVEN_SEGMENT_N_O_0_s1_translator:av_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                                         // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                                           // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                              // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                             // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                              // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                                          // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                              // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                               // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                                // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                                  // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_0_data_master_translator_avalon_universal_master_0_lock;                                                     // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_0_data_master_translator_avalon_universal_master_0_write;                                                    // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_0_data_master_translator_avalon_universal_master_0_read;                                                     // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                                 // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire         cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                              // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                               // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                            // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	wire  [20:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // sram_0_avalon_sram_slave_translator:uav_waitrequest -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_sram_slave_translator:uav_burstcount
	wire  [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_sram_slave_translator:uav_writedata
	wire  [20:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                                   // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_sram_slave_translator:uav_address
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                                     // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_sram_slave_translator:uav_write
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_sram_slave_translator:uav_lock
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_sram_slave_translator:uav_read
	wire  [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // sram_0_avalon_sram_slave_translator:uav_readdata -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // sram_0_avalon_sram_slave_translator:uav_readdatavalid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_sram_slave_translator:uav_debugaccess
	wire   [1:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_sram_slave_translator:uav_byteenable
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                               // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [20:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                            // SWITCH_I_s1_translator:uav_waitrequest -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch_i_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                             // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SWITCH_I_s1_translator:uav_burstcount
	wire  [31:0] switch_i_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                              // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SWITCH_I_s1_translator:uav_writedata
	wire  [20:0] switch_i_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_address -> SWITCH_I_s1_translator:uav_address
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                  // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_write -> SWITCH_I_s1_translator:uav_write
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                   // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SWITCH_I_s1_translator:uav_lock
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                   // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_read -> SWITCH_I_s1_translator:uav_read
	wire  [31:0] switch_i_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                               // SWITCH_I_s1_translator:uav_readdata -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                          // SWITCH_I_s1_translator:uav_readdatavalid -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                            // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SWITCH_I_s1_translator:uav_debugaccess
	wire   [3:0] switch_i_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                             // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SWITCH_I_s1_translator:uav_byteenable
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                     // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                           // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                   // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                            // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                           // SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                  // SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                        // SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                // SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                         // SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                        // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                      // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                       // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                      // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // PUSH_BUTTON_I_s1_translator:uav_waitrequest -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> PUSH_BUTTON_I_s1_translator:uav_burstcount
	wire  [31:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> PUSH_BUTTON_I_s1_translator:uav_writedata
	wire  [20:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_address -> PUSH_BUTTON_I_s1_translator:uav_address
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_write -> PUSH_BUTTON_I_s1_translator:uav_write
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_lock -> PUSH_BUTTON_I_s1_translator:uav_lock
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_read -> PUSH_BUTTON_I_s1_translator:uav_read
	wire  [31:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // PUSH_BUTTON_I_s1_translator:uav_readdata -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // PUSH_BUTTON_I_s1_translator:uav_readdatavalid -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PUSH_BUTTON_I_s1_translator:uav_debugaccess
	wire   [3:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> PUSH_BUTTON_I_s1_translator:uav_byteenable
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // LED_RED_O_s1_translator:uav_waitrequest -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LED_RED_O_s1_translator:uav_burstcount
	wire  [31:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LED_RED_O_s1_translator:uav_writedata
	wire  [20:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_address -> LED_RED_O_s1_translator:uav_address
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_write -> LED_RED_O_s1_translator:uav_write
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LED_RED_O_s1_translator:uav_lock
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_read -> LED_RED_O_s1_translator:uav_read
	wire  [31:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // LED_RED_O_s1_translator:uav_readdata -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // LED_RED_O_s1_translator:uav_readdatavalid -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LED_RED_O_s1_translator:uav_debugaccess
	wire   [3:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LED_RED_O_s1_translator:uav_byteenable
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                         // LED_GREEN_O_s1_translator:uav_waitrequest -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                          // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LED_GREEN_O_s1_translator:uav_burstcount
	wire  [31:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                           // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LED_GREEN_O_s1_translator:uav_writedata
	wire  [20:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_address;                                             // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_address -> LED_GREEN_O_s1_translator:uav_address
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_write;                                               // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_write -> LED_GREEN_O_s1_translator:uav_write
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LED_GREEN_O_s1_translator:uav_lock
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_read -> LED_GREEN_O_s1_translator:uav_read
	wire  [31:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                            // LED_GREEN_O_s1_translator:uav_readdata -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                       // LED_GREEN_O_s1_translator:uav_readdatavalid -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                         // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LED_GREEN_O_s1_translator:uav_debugaccess
	wire   [3:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                          // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LED_GREEN_O_s1_translator:uav_byteenable
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                  // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                        // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                         // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                        // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                               // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                     // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                             // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                      // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                     // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                   // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                    // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                   // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // custom_counter_component_0_avalon_slave_0_translator:uav_waitrequest -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;               // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> custom_counter_component_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> custom_counter_component_0_avalon_slave_0_translator:uav_writedata
	wire  [20:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                  // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> custom_counter_component_0_avalon_slave_0_translator:uav_address
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                    // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> custom_counter_component_0_avalon_slave_0_translator:uav_write
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                     // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> custom_counter_component_0_avalon_slave_0_translator:uav_lock
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                     // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> custom_counter_component_0_avalon_slave_0_translator:uav_read
	wire  [31:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                 // custom_counter_component_0_avalon_slave_0_translator:uav_readdata -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // custom_counter_component_0_avalon_slave_0_translator:uav_readdatavalid -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> custom_counter_component_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;               // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> custom_counter_component_0_avalon_slave_0_translator:uav_byteenable
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;             // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;              // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;             // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // custom_counter_component2_0_avalon_slave_0_translator:uav_waitrequest -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> custom_counter_component2_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> custom_counter_component2_0_avalon_slave_0_translator:uav_writedata
	wire  [20:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> custom_counter_component2_0_avalon_slave_0_translator:uav_address
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> custom_counter_component2_0_avalon_slave_0_translator:uav_write
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> custom_counter_component2_0_avalon_slave_0_translator:uav_lock
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> custom_counter_component2_0_avalon_slave_0_translator:uav_read
	wire  [31:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // custom_counter_component2_0_avalon_slave_0_translator:uav_readdata -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // custom_counter_component2_0_avalon_slave_0_translator:uav_readdatavalid -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> custom_counter_component2_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> custom_counter_component2_0_avalon_slave_0_translator:uav_byteenable
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // SEVEN_SEGMENT_N_O_0_s1_translator:uav_waitrequest -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_burstcount
	wire  [31:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_writedata
	wire  [20:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_address
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_write
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_lock
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_read
	wire  [31:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // SEVEN_SEGMENT_N_O_0_s1_translator:uav_readdata -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // SEVEN_SEGMENT_N_O_0_s1_translator:uav_readdatavalid -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_debugaccess
	wire   [3:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SEVEN_SEGMENT_N_O_0_s1_translator:uav_byteenable
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [93:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                           // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                   // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [93:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                            // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                           // addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                      // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [93:0] cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                       // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                     // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [75:0] sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                                      // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_001:sink_ready -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [93:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                            // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                  // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                          // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [93:0] switch_i_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                   // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         switch_i_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                  // id_router_003:sink_ready -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [93:0] push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_004:sink_ready -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [93:0] led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_005:sink_ready -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                         // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                               // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                       // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [93:0] led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                               // id_router_006:sink_ready -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                    // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [93:0] custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                     // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_007:sink_ready -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [93:0] custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_008:sink_ready -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [93:0] seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_009:sink_ready -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         burst_adapter_source0_endofpacket;                                                                               // burst_adapter:source0_endofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                                     // burst_adapter:source0_valid -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                             // burst_adapter:source0_startofpacket -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] burst_adapter_source0_data;                                                                                      // burst_adapter:source0_data -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                                     // sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [9:0] burst_adapter_source0_channel;                                                                                   // burst_adapter:source0_channel -> sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                                  // rst_controller:reset_out -> [LED_GREEN_O:reset_n, LED_GREEN_O_s1_translator:reset, LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:reset, LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LED_RED_O:reset_n, LED_RED_O_s1_translator:reset, LED_RED_O_s1_translator_avalon_universal_slave_0_agent:reset, LED_RED_O_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PUSH_BUTTON_I:reset_n, PUSH_BUTTON_I_s1_translator:reset, PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:reset, PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SEVEN_SEGMENT_N_O_0:reset_n, SEVEN_SEGMENT_N_O_0_s1_translator:reset, SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:reset, SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SWITCH_I:reset_n, SWITCH_I_s1_translator:reset, SWITCH_I_s1_translator_avalon_universal_slave_0_agent:reset, SWITCH_I_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, custom_counter_component2_0:resetn, custom_counter_component2_0_avalon_slave_0_translator:reset, custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, custom_counter_component_0:resetn, custom_counter_component_0_avalon_slave_0_translator:reset, custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sram_0:reset, sram_0_avalon_sram_slave_translator:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire         cpu_0_jtag_debug_module_reset_reset;                                                                             // cpu_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                                                 // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                       // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                               // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src0_data;                                                                                        // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [9:0] cmd_xbar_demux_src0_channel;                                                                                     // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                                       // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                                 // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                       // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                               // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src1_data;                                                                                        // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [9:0] cmd_xbar_demux_src1_channel;                                                                                     // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                                       // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                             // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                                   // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                           // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src0_data;                                                                                    // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [9:0] cmd_xbar_demux_001_src0_channel;                                                                                 // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                                   // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                             // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                                   // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                           // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src1_data;                                                                                    // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [9:0] cmd_xbar_demux_001_src1_channel;                                                                                 // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                                   // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                             // cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                                   // cmd_xbar_demux_001:src2_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                           // cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src2_data;                                                                                    // cmd_xbar_demux_001:src2_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src2_channel;                                                                                 // cmd_xbar_demux_001:src2_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                             // cmd_xbar_demux_001:src3_endofpacket -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                                   // cmd_xbar_demux_001:src3_valid -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                           // cmd_xbar_demux_001:src3_startofpacket -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src3_data;                                                                                    // cmd_xbar_demux_001:src3_data -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src3_channel;                                                                                 // cmd_xbar_demux_001:src3_channel -> SWITCH_I_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                             // cmd_xbar_demux_001:src4_endofpacket -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                                   // cmd_xbar_demux_001:src4_valid -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                           // cmd_xbar_demux_001:src4_startofpacket -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src4_data;                                                                                    // cmd_xbar_demux_001:src4_data -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src4_channel;                                                                                 // cmd_xbar_demux_001:src4_channel -> PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                             // cmd_xbar_demux_001:src5_endofpacket -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                                   // cmd_xbar_demux_001:src5_valid -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                           // cmd_xbar_demux_001:src5_startofpacket -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src5_data;                                                                                    // cmd_xbar_demux_001:src5_data -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src5_channel;                                                                                 // cmd_xbar_demux_001:src5_channel -> LED_RED_O_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                             // cmd_xbar_demux_001:src6_endofpacket -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                                   // cmd_xbar_demux_001:src6_valid -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                           // cmd_xbar_demux_001:src6_startofpacket -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src6_data;                                                                                    // cmd_xbar_demux_001:src6_data -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src6_channel;                                                                                 // cmd_xbar_demux_001:src6_channel -> LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                             // cmd_xbar_demux_001:src7_endofpacket -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                                   // cmd_xbar_demux_001:src7_valid -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                           // cmd_xbar_demux_001:src7_startofpacket -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src7_data;                                                                                    // cmd_xbar_demux_001:src7_data -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src7_channel;                                                                                 // cmd_xbar_demux_001:src7_channel -> custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                             // cmd_xbar_demux_001:src8_endofpacket -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                                   // cmd_xbar_demux_001:src8_valid -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                           // cmd_xbar_demux_001:src8_startofpacket -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src8_data;                                                                                    // cmd_xbar_demux_001:src8_data -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src8_channel;                                                                                 // cmd_xbar_demux_001:src8_channel -> custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                             // cmd_xbar_demux_001:src9_endofpacket -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                                   // cmd_xbar_demux_001:src9_valid -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                                           // cmd_xbar_demux_001:src9_startofpacket -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src9_data;                                                                                    // cmd_xbar_demux_001:src9_data -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_demux_001_src9_channel;                                                                                 // cmd_xbar_demux_001:src9_channel -> SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                                 // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                       // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                               // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [93:0] rsp_xbar_demux_src0_data;                                                                                        // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [9:0] rsp_xbar_demux_src0_channel;                                                                                     // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                       // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                                 // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                                       // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                               // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [93:0] rsp_xbar_demux_src1_data;                                                                                        // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [9:0] rsp_xbar_demux_src1_channel;                                                                                     // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                                       // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                             // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                                   // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                           // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [93:0] rsp_xbar_demux_001_src0_data;                                                                                    // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [9:0] rsp_xbar_demux_001_src0_channel;                                                                                 // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                                   // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                             // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                                   // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                           // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [93:0] rsp_xbar_demux_001_src1_data;                                                                                    // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [9:0] rsp_xbar_demux_001_src1_channel;                                                                                 // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                                   // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                             // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                                   // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                           // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [93:0] rsp_xbar_demux_002_src0_data;                                                                                    // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [9:0] rsp_xbar_demux_002_src0_channel;                                                                                 // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                                   // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                             // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                                   // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                           // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [93:0] rsp_xbar_demux_003_src0_data;                                                                                    // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [9:0] rsp_xbar_demux_003_src0_channel;                                                                                 // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                                   // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                             // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                                   // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                           // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [93:0] rsp_xbar_demux_004_src0_data;                                                                                    // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [9:0] rsp_xbar_demux_004_src0_channel;                                                                                 // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                                   // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                             // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                                   // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                           // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [93:0] rsp_xbar_demux_005_src0_data;                                                                                    // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [9:0] rsp_xbar_demux_005_src0_channel;                                                                                 // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                                   // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                             // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                                   // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                           // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [93:0] rsp_xbar_demux_006_src0_data;                                                                                    // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [9:0] rsp_xbar_demux_006_src0_channel;                                                                                 // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                                   // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                             // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                                   // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                           // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [93:0] rsp_xbar_demux_007_src0_data;                                                                                    // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [9:0] rsp_xbar_demux_007_src0_channel;                                                                                 // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                                   // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                             // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                                   // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                           // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [93:0] rsp_xbar_demux_008_src0_data;                                                                                    // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [9:0] rsp_xbar_demux_008_src0_channel;                                                                                 // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                                   // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                             // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                                   // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                                           // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [93:0] rsp_xbar_demux_009_src0_data;                                                                                    // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [9:0] rsp_xbar_demux_009_src0_channel;                                                                                 // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                                   // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         addr_router_src_endofpacket;                                                                                     // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                                           // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                                   // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [93:0] addr_router_src_data;                                                                                            // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [9:0] addr_router_src_channel;                                                                                         // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                                           // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                                    // rsp_xbar_mux:src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                          // rsp_xbar_mux:src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                                  // rsp_xbar_mux:src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [93:0] rsp_xbar_mux_src_data;                                                                                           // rsp_xbar_mux:src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [9:0] rsp_xbar_mux_src_channel;                                                                                        // rsp_xbar_mux:src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                                          // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                                 // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                                       // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                               // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [93:0] addr_router_001_src_data;                                                                                        // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [9:0] addr_router_001_src_channel;                                                                                     // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                                       // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                                // rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                                      // rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                              // rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [93:0] rsp_xbar_mux_001_src_data;                                                                                       // rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [9:0] rsp_xbar_mux_001_src_channel;                                                                                    // rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                                      // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                                    // cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                          // cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                                  // cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_src_data;                                                                                           // cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [9:0] cmd_xbar_mux_src_channel;                                                                                        // cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                          // cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                                       // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                             // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                                     // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [93:0] id_router_src_data;                                                                                              // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [9:0] id_router_src_channel;                                                                                           // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                             // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_001_src2_ready;                                                                                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire         id_router_002_src_endofpacket;                                                                                   // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                         // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                                 // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [93:0] id_router_002_src_data;                                                                                          // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [9:0] id_router_002_src_channel;                                                                                       // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                         // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                                   // SWITCH_I_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                                   // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                         // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                                 // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [93:0] id_router_003_src_data;                                                                                          // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [9:0] id_router_003_src_channel;                                                                                       // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                         // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                                   // PUSH_BUTTON_I_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                                   // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                         // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                                 // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [93:0] id_router_004_src_data;                                                                                          // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [9:0] id_router_004_src_channel;                                                                                       // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                         // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                                   // LED_RED_O_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                                   // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                         // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                                 // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [93:0] id_router_005_src_data;                                                                                          // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [9:0] id_router_005_src_channel;                                                                                       // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                         // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                                   // LED_GREEN_O_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                                   // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                         // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                                 // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [93:0] id_router_006_src_data;                                                                                          // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [9:0] id_router_006_src_channel;                                                                                       // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                         // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                                   // custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                                   // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                         // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                                 // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [93:0] id_router_007_src_data;                                                                                          // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [9:0] id_router_007_src_channel;                                                                                       // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                         // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                                   // custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                                   // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                         // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                                 // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [93:0] id_router_008_src_data;                                                                                          // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [9:0] id_router_008_src_channel;                                                                                       // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                         // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                                   // SEVEN_SEGMENT_N_O_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                                   // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                                         // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                                 // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [93:0] id_router_009_src_data;                                                                                          // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [9:0] id_router_009_src_channel;                                                                                       // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                                         // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                                // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                                      // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                              // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [93:0] cmd_xbar_mux_001_src_data;                                                                                       // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [9:0] cmd_xbar_mux_001_src_channel;                                                                                    // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                                      // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire         width_adapter_src_endofpacket;                                                                                   // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                                         // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                                 // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [75:0] width_adapter_src_data;                                                                                          // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                                         // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [9:0] width_adapter_src_channel;                                                                                       // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_001_src_endofpacket;                                                                                   // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_001_src_valid;                                                                                         // id_router_001:src_valid -> width_adapter_001:in_valid
	wire         id_router_001_src_startofpacket;                                                                                 // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [75:0] id_router_001_src_data;                                                                                          // id_router_001:src_data -> width_adapter_001:in_data
	wire   [9:0] id_router_001_src_channel;                                                                                       // id_router_001:src_channel -> width_adapter_001:in_channel
	wire         id_router_001_src_ready;                                                                                         // width_adapter_001:in_ready -> id_router_001:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                               // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                                     // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                             // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [93:0] width_adapter_001_src_data;                                                                                      // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire         width_adapter_001_src_ready;                                                                                     // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [9:0] width_adapter_001_src_channel;                                                                                   // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire         irq_mapper_receiver0_irq;                                                                                        // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                                        // PUSH_BUTTON_I:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                                        // custom_counter_component_0:counter_expire_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                                        // custom_counter_component2_0:counter_expire_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                                        // SWITCH_I:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_0_d_irq_irq;                                                                                                 // irq_mapper:sender_irq -> cpu_0:d_irq

	experiment1b_sram_0 sram_0 (
		.clk           (clk_50_i_in_clk),                                                       //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                        //  clock_reset_reset.reset
		.SRAM_DQ       (sram_0_external_interface_DQ),                                          // external_interface.export
		.SRAM_ADDR     (sram_0_external_interface_ADDR),                                        //                   .export
		.SRAM_LB_N     (sram_0_external_interface_LB_N),                                        //                   .export
		.SRAM_UB_N     (sram_0_external_interface_UB_N),                                        //                   .export
		.SRAM_CE_N     (sram_0_external_interface_CE_N),                                        //                   .export
		.SRAM_OE_N     (sram_0_external_interface_OE_N),                                        //                   .export
		.SRAM_WE_N     (sram_0_external_interface_WE_N),                                        //                   .export
		.address       (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	experiment1b_cpu_0 cpu_0 (
		.clk                                   (clk_50_i_in_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (cpu_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.d_irq                                 (cpu_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	experiment1b_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_50_i_in_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	experiment1b_SWITCH_I switch_i (
		.clk        (clk_50_i_in_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (switch_i_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch_i_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch_i_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch_i_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch_i_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch_i_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                               //                 irq.irq
	);

	experiment1b_PUSH_BUTTON_I push_button_i (
		.clk        (clk_50_i_in_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (push_button_i_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~push_button_i_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (push_button_i_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (push_button_i_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (push_button_i_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (push_button_i_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                                    //                 irq.irq
	);

	experiment1b_LED_RED_O led_red_o (
		.clk        (clk_50_i_in_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (led_red_o_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_red_o_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_red_o_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_red_o_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_red_o_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_red_o_external_connection_export)                    // external_connection.export
	);

	experiment1b_LED_GREEN_O led_green_o (
		.clk        (clk_50_i_in_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (led_green_o_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_green_o_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_green_o_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_green_o_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_green_o_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_green_o_external_connection_export)                    // external_connection.export
	);

	custom_counter_component custom_counter_component_0 (
		.address            (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //   avalon_slave_0.address
		.chipselect         (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.read               (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                 .read
		.write              (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                 .write
		.readdata           (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.writedata          (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.clock              (clk_50_i_in_clk),                                                                     //       clock_sink.clk
		.resetn             (~rst_controller_reset_out_reset),                                                     //       reset_sink.reset_n
		.counter_expire_irq (irq_mapper_receiver2_irq)                                                             // interrupt_sender.irq
	);

	custom_counter_component custom_counter_component2_0 (
		.address            (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //   avalon_slave_0.address
		.chipselect         (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.read               (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                 .read
		.write              (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                 .write
		.readdata           (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.writedata          (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.clock              (clk_50_i_in_clk),                                                                      //       clock_sink.clk
		.resetn             (~rst_controller_reset_out_reset),                                                      //       reset_sink.reset_n
		.counter_expire_irq (irq_mapper_receiver3_irq)                                                              // interrupt_sender.irq
	);

	experiment1b_SEVEN_SEGMENT_N_O_0 seven_segment_n_o_0 (
		.clk        (clk_50_i_in_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                  //               reset.reset_n
		.address    (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (seven_segment_n_o_0_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                   (clk_50_i_in_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_readdatavalid      (),                                                                            //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_0_data_master_translator (
		.clk                   (clk_50_i_in_clk),                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_0_data_master_read),                                               //                          .read
		.av_readdata           (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_0_data_master_write),                                              //                          .write
		.av_writedata          (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_0_jtag_debug_module_translator (
		.clk                   (clk_50_i_in_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_0_avalon_sram_slave_translator (
		.clk                   (clk_50_i_in_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sram_0_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clk_50_i_in_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_i_s1_translator (
		.clk                   (clk_50_i_in_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_i_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (switch_i_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (switch_i_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (switch_i_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (switch_i_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) push_button_i_s1_translator (
		.clk                   (clk_50_i_in_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (push_button_i_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (push_button_i_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (push_button_i_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (push_button_i_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (push_button_i_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_red_o_s1_translator (
		.clk                   (clk_50_i_in_clk),                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_red_o_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_red_o_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_red_o_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_red_o_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_red_o_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_green_o_s1_translator (
		.clk                   (clk_50_i_in_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address           (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_green_o_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_green_o_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_green_o_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_green_o_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_green_o_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) custom_counter_component_0_avalon_slave_0_translator (
		.clk                   (clk_50_i_in_clk),                                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                       //                    reset.reset
		.uav_address           (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (custom_counter_component_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                                     //              (terminated)
		.av_lock               (),                                                                                                     //              (terminated)
		.av_clken              (),                                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) custom_counter_component2_0_avalon_slave_0_translator (
		.clk                   (clk_50_i_in_clk),                                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                        //                    reset.reset
		.uav_address           (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (custom_counter_component2_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                                      //              (terminated)
		.av_lock               (),                                                                                                      //              (terminated)
		.av_clken              (),                                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seven_segment_n_o_0_s1_translator (
		.clk                   (clk_50_i_in_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (seven_segment_n_o_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                  //              (terminated)
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (75),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_50_i_in_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (75),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (10),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_50_i_in_clk),                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (57),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (38),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (39),
		.PKT_TRANS_POSTED          (40),
		.PKT_TRANS_WRITE           (41),
		.PKT_TRANS_READ            (42),
		.PKT_TRANS_LOCK            (43),
		.PKT_SRC_ID_H              (61),
		.PKT_SRC_ID_L              (58),
		.PKT_DEST_ID_H             (65),
		.PKT_DEST_ID_L             (62),
		.PKT_BURSTWRAP_H           (50),
		.PKT_BURSTWRAP_L           (48),
		.PKT_BYTE_CNT_H            (47),
		.PKT_BYTE_CNT_L            (45),
		.PKT_PROTECTION_H          (69),
		.PKT_PROTECTION_L          (67),
		.PKT_RESPONSE_STATUS_H     (75),
		.PKT_RESPONSE_STATUS_L     (74),
		.PKT_BURST_SIZE_H          (53),
		.PKT_BURST_SIZE_L          (51),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                 //                .channel
		.rf_sink_ready           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_i_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_i_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                  //                .channel
		.rf_sink_ready           (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_i_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) push_button_i_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (push_button_i_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                       //                .channel
		.rf_sink_ready           (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (push_button_i_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (push_button_i_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (push_button_i_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_red_o_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_red_o_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                   //                .channel
		.rf_sink_ready           (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_red_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_red_o_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_red_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_green_o_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_green_o_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                     //                .channel
		.rf_sink_ready           (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_green_o_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_green_o_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_green_o_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                 //       clk_reset.reset
		.m0_address              (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                                //                .channel
		.rf_sink_ready           (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                 // clk_reset.reset
		.in_data           (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                                           // (terminated)
		.csr_readdata      (),                                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                           // (terminated)
		.almost_full_data  (),                                                                                                               // (terminated)
		.almost_empty_data (),                                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                                           // (terminated)
		.out_empty         (),                                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                                           // (terminated)
		.out_error         (),                                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                                           // (terminated)
		.out_channel       ()                                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                  //       clk_reset.reset
		.m0_address              (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                                 //                .channel
		.rf_sink_ready           (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                  // clk_reset.reset
		.in_data           (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                            // (terminated)
		.almost_full_data  (),                                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                                            // (terminated)
		.out_empty         (),                                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                                            // (terminated)
		.out_error         (),                                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                                            // (terminated)
		.out_channel       ()                                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (79),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (80),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (10),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_50_i_in_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                             //                .channel
		.rf_sink_ready           (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_50_i_in_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	experiment1b_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	experiment1b_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	experiment1b_id_router id_router (
		.sink_ready         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	experiment1b_id_router_001 id_router_001 (
		.sink_ready         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_0_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                             //       src.ready
		.src_valid          (id_router_001_src_valid),                                                             //          .valid
		.src_data           (id_router_001_src_data),                                                              //          .data
		.src_channel        (id_router_001_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                        //          .endofpacket
	);

	experiment1b_id_router_002 id_router_002 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                             //          .endofpacket
	);

	experiment1b_id_router_002 id_router_003 (
		.sink_ready         (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_i_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                //          .valid
		.src_data           (id_router_003_src_data),                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                           //          .endofpacket
	);

	experiment1b_id_router_002 id_router_004 (
		.sink_ready         (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (push_button_i_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                     //       src.ready
		.src_valid          (id_router_004_src_valid),                                                     //          .valid
		.src_data           (id_router_004_src_data),                                                      //          .data
		.src_channel        (id_router_004_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                //          .endofpacket
	);

	experiment1b_id_router_002 id_router_005 (
		.sink_ready         (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_red_o_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                 //       src.ready
		.src_valid          (id_router_005_src_valid),                                                 //          .valid
		.src_data           (id_router_005_src_data),                                                  //          .data
		.src_channel        (id_router_005_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                            //          .endofpacket
	);

	experiment1b_id_router_002 id_router_006 (
		.sink_ready         (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_green_o_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                   //       src.ready
		.src_valid          (id_router_006_src_valid),                                                   //          .valid
		.src_data           (id_router_006_src_data),                                                    //          .data
		.src_channel        (id_router_006_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                              //          .endofpacket
	);

	experiment1b_id_router_002 id_router_007 (
		.sink_ready         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (custom_counter_component_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                              //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                              //          .valid
		.src_data           (id_router_007_src_data),                                                                               //          .data
		.src_channel        (id_router_007_src_channel),                                                                            //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                                      //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                                         //          .endofpacket
	);

	experiment1b_id_router_002 id_router_008 (
		.sink_ready         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (custom_counter_component2_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                               //          .valid
		.src_data           (id_router_008_src_data),                                                                                //          .data
		.src_channel        (id_router_008_src_channel),                                                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                          //          .endofpacket
	);

	experiment1b_id_router_002 id_router_009 (
		.sink_ready         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seven_segment_n_o_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_50_i_in_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                           //       src.ready
		.src_valid          (id_router_009_src_valid),                                                           //          .valid
		.src_data           (id_router_009_src_data),                                                            //          .data
		.src_channel        (id_router_009_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                      //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (38),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (57),
		.PKT_BYTE_CNT_H            (47),
		.PKT_BYTE_CNT_L            (45),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (53),
		.PKT_BURST_SIZE_L          (51),
		.PKT_BURST_TYPE_H          (55),
		.PKT_BURST_TYPE_L          (54),
		.PKT_BURSTWRAP_H           (50),
		.PKT_BURSTWRAP_L           (48),
		.PKT_TRANS_COMPRESSED_READ (39),
		.PKT_TRANS_WRITE           (41),
		.PKT_TRANS_READ            (42),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (10),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (50),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk_50_i_in_clk),                     //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~clk_50_i_in_reset_reset_n),          // reset_in0.reset
		.reset_in1  (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_50_i_in_clk),                     //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	experiment1b_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_50_i_in_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	experiment1b_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //      src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //      src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.src8_ready         (cmd_xbar_demux_001_src8_ready),         //      src8.ready
		.src8_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.src8_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.src8_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.src8_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.src8_endofpacket   (cmd_xbar_demux_001_src8_endofpacket),   //          .endofpacket
		.src9_ready         (cmd_xbar_demux_001_src9_ready),         //      src9.ready
		.src9_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.src9_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.src9_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.src9_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.src9_endofpacket   (cmd_xbar_demux_001_src9_endofpacket)    //          .endofpacket
	);

	experiment1b_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_50_i_in_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_50_i_in_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	experiment1b_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clk_50_i_in_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	experiment1b_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (clk_50_i_in_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_50_i_in_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	experiment1b_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_50_i_in_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready         (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready         (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (56),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (65),
		.IN_PKT_BYTE_CNT_L             (63),
		.IN_PKT_TRANS_COMPRESSED_READ  (57),
		.IN_PKT_BURSTWRAP_H            (68),
		.IN_PKT_BURSTWRAP_L            (66),
		.IN_PKT_BURST_SIZE_H           (71),
		.IN_PKT_BURST_SIZE_L           (69),
		.IN_PKT_RESPONSE_STATUS_H      (93),
		.IN_PKT_RESPONSE_STATUS_L      (92),
		.IN_PKT_TRANS_EXCLUSIVE        (62),
		.IN_PKT_BURST_TYPE_H           (73),
		.IN_PKT_BURST_TYPE_L           (72),
		.IN_ST_DATA_W                  (94),
		.OUT_PKT_ADDR_H                (38),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (47),
		.OUT_PKT_BYTE_CNT_L            (45),
		.OUT_PKT_TRANS_COMPRESSED_READ (39),
		.OUT_PKT_BURST_SIZE_H          (53),
		.OUT_PKT_BURST_SIZE_L          (51),
		.OUT_PKT_RESPONSE_STATUS_H     (75),
		.OUT_PKT_RESPONSE_STATUS_L     (74),
		.OUT_PKT_TRANS_EXCLUSIVE       (44),
		.OUT_PKT_BURST_TYPE_H          (55),
		.OUT_PKT_BURST_TYPE_L          (54),
		.OUT_ST_DATA_W                 (76),
		.ST_CHANNEL_W                  (10),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clk_50_i_in_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (38),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (47),
		.IN_PKT_BYTE_CNT_L             (45),
		.IN_PKT_TRANS_COMPRESSED_READ  (39),
		.IN_PKT_BURSTWRAP_H            (50),
		.IN_PKT_BURSTWRAP_L            (48),
		.IN_PKT_BURST_SIZE_H           (53),
		.IN_PKT_BURST_SIZE_L           (51),
		.IN_PKT_RESPONSE_STATUS_H      (75),
		.IN_PKT_RESPONSE_STATUS_L      (74),
		.IN_PKT_TRANS_EXCLUSIVE        (44),
		.IN_PKT_BURST_TYPE_H           (55),
		.IN_PKT_BURST_TYPE_L           (54),
		.IN_ST_DATA_W                  (76),
		.OUT_PKT_ADDR_H                (56),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (65),
		.OUT_PKT_BYTE_CNT_L            (63),
		.OUT_PKT_TRANS_COMPRESSED_READ (57),
		.OUT_PKT_BURST_SIZE_H          (71),
		.OUT_PKT_BURST_SIZE_L          (69),
		.OUT_PKT_RESPONSE_STATUS_H     (93),
		.OUT_PKT_RESPONSE_STATUS_L     (92),
		.OUT_PKT_TRANS_EXCLUSIVE       (62),
		.OUT_PKT_BURST_TYPE_H          (73),
		.OUT_PKT_BURST_TYPE_L          (72),
		.OUT_ST_DATA_W                 (94),
		.ST_CHANNEL_W                  (10),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (clk_50_i_in_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	experiment1b_irq_mapper irq_mapper (
		.clk           (clk_50_i_in_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

endmodule
